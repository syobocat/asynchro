module main

import service.database

fn init_db() ! {
	println('Initializing the database...')
	database.init_db()!
	println('Database initialized.')
}
